module tetromino_rom ( input [6:0]	addr,
						output [3:0]	data
					 );

	parameter ADDR_WIDTH = 7;
   parameter DATA_WIDTH =  4;
	logic [ADDR_WIDTH-1:0] addr_reg;
	
	// Orientations, addr[1:0]:
	// 00: Upright
	// 01: Turned right clockwise
	// 10: Upside down
	// 11: Turned left counterclockwise
	
	//Blocks
	// 000: I
	// 001: Left-L
	// 010: Right-L
	// 011: Block
	// 100: S
	// 101: T
	// 110: Z
	
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		//I
		//00
		4'b0000,
		4'b0000,
		4'b1111,
		4'b0000,
		//01
		4'b0010,
		4'b0010,
		4'b0010,
		4'b0010,
		//10
		4'b0000,
		4'b0000,
		4'b1111,
		4'b0000,
		//11
		4'b0010,
		4'b0010,
		4'b0010,
		4'b0010,
		//Left-L
		//00
		4'b0000,
		4'b1000,
		4'b1110,
		4'b0000,
		//01
		4'b1100,
		4'b1000,
		4'b1000,
		4'b0000,
		//10
		4'b0000,
		4'b1110,
		4'b0010,
		4'b0000,
		//11
		4'b0100,
		4'b0100,
		4'b1100,
		4'b0000,
		//Right-L
		//00
		4'b0000,
		4'b0010,
		4'b1110,
		4'b0000,
		//01
		4'b0100,
		4'b0100,
		4'b0110,
		4'b0000,
		//10
		4'b0000,
		4'b1110,
		4'b1000,
		4'b0000,
		//11
		4'b0110,
		4'b0010,
		4'b0010,
		4'b0000,
		//Block
		//00
		4'b0000,
		4'b0110,
		4'b0110,
		4'b0000,
		//01
		4'b0000,
		4'b0110,
		4'b0110,
		4'b0000,
		//10
		4'b0000,
		4'b0110,
		4'b0110,
		4'b0000,
		//11
		4'b0000,
		4'b0110,
		4'b0110,
		4'b0000,
		//S
		//00
		4'b0000,
		4'b0110,
		4'b1100,
		4'b0000,
		//01
		4'b0000,
		4'b0100,
		4'b0110,
		4'b0010,
		//10
		4'b0000,
		4'b0110,
		4'b1100,
		4'b0000,
		//11
		4'b0000,
		4'b0100,
		4'b0110,
		4'b0010,
		//T
		//00
		4'b0000,
		4'b0100,
		4'b1110,
		4'b0000,
		//01
		4'b0000,
		4'b0100,
		4'b0110,
		4'b0100,
		//10
		4'b0000,
		4'b1110,
		4'b0100,
		4'b0000,
		//11
		4'b0000,
		4'b0100,
		4'b1100,
		4'b0100,
		//Z
		//00
		4'b0000,
		4'b1100,
		4'b0110,
		4'b0000,
		//01
		4'b0000,
		4'b0010,
		4'b0110,
		4'b0100,
		//10
		4'b0000,
		4'b1100,
		4'b0110,
		4'b0000,
		//11
		4'b0000,
		4'b0010,
		4'b0110,
		4'b0100,
		//I
		//00
		4'b0000,
		4'b0000,
		4'b1111,
		4'b0000,
		//01
		4'b0010,
		4'b0010,
		4'b0010,
		4'b0010,
		//10
		4'b0000,
		4'b0000,
		4'b1111,
		4'b0000,
		//11
		4'b0010,
		4'b0010,
		4'b0010,
		4'b0010
	};
	
	assign data = ROM[addr];
	
endmodule